library verilog;
use verilog.vl_types.all;
entity sramif_vlg_vec_tst is
end sramif_vlg_vec_tst;
